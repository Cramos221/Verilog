


package test_pkg;

  

  
  `include "uvm_macros.svh"
  `include "interface.svh"
  `include "sequence_item.svh"
  `include "sequencer.svh"
  `include "sequence.svh"
  `include "driver.svh"
  `include "monitor.svh"
  `include "agent.svh"
  `include "env.svh"
  `include "test.svh"
  `include "scoreboard.svh"
 

endpackage
  
