interface seq_if;
  
  
   logic in;
  logic clk;
  logic reset;
  logic out;

endinterface