// A coleção de portas de sinal para DUT e testbench
interface our_interface (input logic clk); 
  
 
  logic [7:0] input_1;
  logic [7:0] input_2;
  logic [7:0] input_3;
  logic [7:0] input_4;
  logic [7:0] input_5;
  logic [7:0] input_6;
  logic [7:0] input_7;
  logic [7:0] input_8;
  
  logic [7:0] out1;
  logic [7:0] out2;
  logic [7:0] out3;
  logic [7:0] out4;
  logic [7:0] out5;
  logic [7:0] out6;
  logic [7:0] out7;
  logic [7:0] out8;
  
  
endinterface: our_interface

